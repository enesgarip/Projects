module br_j_control(branch,status,out_j_control);
input [1:0] branch,status;
output out_j_control;
reg[1:0] out_j_control;
reg clk;
initial
begin
clk = 0;
forever #20  clk=~clk;
end

always @(posedge clk)
begin
if((~branch[1]) & (~branch[0])) out_j_control=2'b00;					//Jump instructionlar? i�in kosulsuz atlama
else if(branch[1] & branch[0]&status[1] & (~status[0])) out_j_control=2'b11;		// beq i�in atlama
else if(branch[1] & (~branch[0]) & (~status[0])) out_j_control=2'b11;			// bgez i�in atlama
else if((~branch[0]) & branch[1] & status[1]) out_j_control=2'b10;			// balz i�in atlama
else out_j_control=2'b00;
end

endmodule

/*
	00 - Ordinar path
	01 - Jumpaddress ( 26 bit )
	10 - Balz ( 26 bit ) 
	11 - brench pc-relative

*/
